module tb_sample_test;

    initial
    begin
        $display("Test has been run!");
        $finish();
    end

endmodule

