// Module takes in data from a full block of registers. Selects the correct
// elements from this block based on vsew and address.

module element_selector (
    output logic [127:0] data_out,
    input wire [127:0] block_data,
    input wire [4:0] addr,
    input wire [1:0] vsew
);



endmodule
